module out_port_seg(in,out1,out0);
	input 	[31: 0] in				;
	output 	[ 6: 0] out1,out0		;
	
	reg 		[ 3: 0] num5,num4,num3,num2,num1,num0;

	sevenseg display_1( num1, out1 );
	sevenseg display_0( num0, out0 );
	
	always @ (in)
	begin
		num1 = ( in / 10 ) % 10;
		num0 = in % 10;
	end
	
endmodule

module sevenseg(data, ledsegments);
	input 	[ 3: 0] 		data				;
	output 					ledsegments		;
	reg 		[ 6: 0] 		ledsegments		;
	
	always @ (*)
		case(data)
			0: ledsegments = 7'b100_0000;
			1: ledsegments = 7'b111_1001;
			2: ledsegments = 7'b010_0100;
			3: ledsegments = 7'b011_0000;
			4: ledsegments = 7'b001_1001;
			5: ledsegments = 7'b001_0010;
			6: ledsegments = 7'b000_0010;
			7: ledsegments = 7'b111_1000;
			8: ledsegments = 7'b000_0000;
			9: ledsegments = 7'b001_0000;
			default: ledsegments = 7'b111_1111;
		endcase
endmodule